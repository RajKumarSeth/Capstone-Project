module add_sub(a,b,c,sum,carry);
parameter n=8;
input [n-1:0] a,b;
input c;
output [n-1:0] sum;
output carry;
wire [n-2:0] co;
wire [n-1:0] x;
xor xor0(x[0],b[0],c);
xor xor1(x[1],b[1],c);
xor xor2(x[2],b[2],c);
xor xor3(x[3],b[3],c);
xor xor4(x[4],b[4],c);
xor xor5(x[5],b[5],c);
xor xor6(x[6],b[6],c);
xor xor7(x[7],b[7],c);
full_adder fa0(.a(a[0]),.b(x[0]),.c(c),.sum(sum[0]),.carry(co[0]));
full_adder fa1(.a(a[1]),.b(x[1]),.c(co[0]),.sum(sum[1]),.carry(co[1]));
full_adder fa2(.a(a[2]),.b(x[2]),.c(co[1]),.sum(sum[2]),.carry(co[2]));
full_adder fa3(.a(a[3]),.b(x[3]),.c(co[2]),.sum(sum[3]),.carry(co[3]));
full_adder fa4(.a(a[4]),.b(x[4]),.c(co[3]),.sum(sum[4]),.carry(co[4]));
full_adder fa5(.a(a[5]),.b(x[5]),.c(co[4]),.sum(sum[5]),.carry(co[5]));
full_adder fa6(.a(a[6]),.b(x[6]),.c(co[5]),.sum(sum[6]),.carry(co[6]));
full_adder fa7(.a(a[7]),.b(x[7]),.c(co[6]),.sum(sum[7]),.carry(carry));
endmodule
